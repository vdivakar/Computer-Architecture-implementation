module first;
  initial
  begin 
    $display("hello");
  end
endmodule
